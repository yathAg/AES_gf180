magic
tech gf180mcuD
magscale 1 5
timestamp 1701671474
<< obsm1 >>
rect 672 855 259280 278350
<< metal2 >>
rect 12320 0 12376 400
rect 13104 0 13160 400
rect 13888 0 13944 400
rect 14672 0 14728 400
rect 15456 0 15512 400
rect 16240 0 16296 400
rect 17024 0 17080 400
rect 17808 0 17864 400
rect 18592 0 18648 400
rect 19376 0 19432 400
rect 20160 0 20216 400
rect 20944 0 21000 400
rect 21728 0 21784 400
rect 22512 0 22568 400
rect 23296 0 23352 400
rect 24080 0 24136 400
rect 24864 0 24920 400
rect 25648 0 25704 400
rect 26432 0 26488 400
rect 27216 0 27272 400
rect 28000 0 28056 400
rect 28784 0 28840 400
rect 29568 0 29624 400
rect 30352 0 30408 400
rect 31136 0 31192 400
rect 31920 0 31976 400
rect 32704 0 32760 400
rect 33488 0 33544 400
rect 34272 0 34328 400
rect 35056 0 35112 400
rect 35840 0 35896 400
rect 36624 0 36680 400
rect 37408 0 37464 400
rect 38192 0 38248 400
rect 38976 0 39032 400
rect 39760 0 39816 400
rect 40544 0 40600 400
rect 41328 0 41384 400
rect 42112 0 42168 400
rect 42896 0 42952 400
rect 43680 0 43736 400
rect 44464 0 44520 400
rect 45248 0 45304 400
rect 46032 0 46088 400
rect 46816 0 46872 400
rect 47600 0 47656 400
rect 48384 0 48440 400
rect 49168 0 49224 400
rect 49952 0 50008 400
rect 50736 0 50792 400
rect 51520 0 51576 400
rect 52304 0 52360 400
rect 53088 0 53144 400
rect 53872 0 53928 400
rect 54656 0 54712 400
rect 55440 0 55496 400
rect 56224 0 56280 400
rect 57008 0 57064 400
rect 57792 0 57848 400
rect 58576 0 58632 400
rect 59360 0 59416 400
rect 60144 0 60200 400
rect 60928 0 60984 400
rect 61712 0 61768 400
rect 62496 0 62552 400
rect 63280 0 63336 400
rect 64064 0 64120 400
rect 64848 0 64904 400
rect 65632 0 65688 400
rect 66416 0 66472 400
rect 67200 0 67256 400
rect 67984 0 68040 400
rect 68768 0 68824 400
rect 69552 0 69608 400
rect 70336 0 70392 400
rect 71120 0 71176 400
rect 71904 0 71960 400
rect 72688 0 72744 400
rect 73472 0 73528 400
rect 74256 0 74312 400
rect 75040 0 75096 400
rect 75824 0 75880 400
rect 76608 0 76664 400
rect 77392 0 77448 400
rect 78176 0 78232 400
rect 78960 0 79016 400
rect 79744 0 79800 400
rect 80528 0 80584 400
rect 81312 0 81368 400
rect 82096 0 82152 400
rect 82880 0 82936 400
rect 83664 0 83720 400
rect 84448 0 84504 400
rect 85232 0 85288 400
rect 86016 0 86072 400
rect 86800 0 86856 400
rect 87584 0 87640 400
rect 88368 0 88424 400
rect 89152 0 89208 400
rect 89936 0 89992 400
rect 90720 0 90776 400
rect 91504 0 91560 400
rect 92288 0 92344 400
rect 93072 0 93128 400
rect 93856 0 93912 400
rect 94640 0 94696 400
rect 95424 0 95480 400
rect 96208 0 96264 400
rect 96992 0 97048 400
rect 97776 0 97832 400
rect 98560 0 98616 400
rect 99344 0 99400 400
rect 100128 0 100184 400
rect 100912 0 100968 400
rect 101696 0 101752 400
rect 102480 0 102536 400
rect 103264 0 103320 400
rect 104048 0 104104 400
rect 104832 0 104888 400
rect 105616 0 105672 400
rect 106400 0 106456 400
rect 107184 0 107240 400
rect 107968 0 108024 400
rect 108752 0 108808 400
rect 109536 0 109592 400
rect 110320 0 110376 400
rect 111104 0 111160 400
rect 111888 0 111944 400
rect 112672 0 112728 400
rect 113456 0 113512 400
rect 114240 0 114296 400
rect 115024 0 115080 400
rect 115808 0 115864 400
rect 116592 0 116648 400
rect 117376 0 117432 400
rect 118160 0 118216 400
rect 118944 0 119000 400
rect 119728 0 119784 400
rect 120512 0 120568 400
rect 121296 0 121352 400
rect 122080 0 122136 400
rect 122864 0 122920 400
rect 123648 0 123704 400
rect 124432 0 124488 400
rect 125216 0 125272 400
rect 126000 0 126056 400
rect 126784 0 126840 400
rect 127568 0 127624 400
rect 128352 0 128408 400
rect 129136 0 129192 400
rect 129920 0 129976 400
rect 130704 0 130760 400
rect 131488 0 131544 400
rect 132272 0 132328 400
rect 133056 0 133112 400
rect 133840 0 133896 400
rect 134624 0 134680 400
rect 135408 0 135464 400
rect 136192 0 136248 400
rect 136976 0 137032 400
rect 137760 0 137816 400
rect 138544 0 138600 400
rect 139328 0 139384 400
rect 140112 0 140168 400
rect 140896 0 140952 400
rect 141680 0 141736 400
rect 142464 0 142520 400
rect 143248 0 143304 400
rect 144032 0 144088 400
rect 144816 0 144872 400
rect 145600 0 145656 400
rect 146384 0 146440 400
rect 147168 0 147224 400
rect 147952 0 148008 400
rect 148736 0 148792 400
rect 149520 0 149576 400
rect 150304 0 150360 400
rect 151088 0 151144 400
rect 151872 0 151928 400
rect 152656 0 152712 400
rect 153440 0 153496 400
rect 154224 0 154280 400
rect 155008 0 155064 400
rect 155792 0 155848 400
rect 156576 0 156632 400
rect 157360 0 157416 400
rect 158144 0 158200 400
rect 158928 0 158984 400
rect 159712 0 159768 400
rect 160496 0 160552 400
rect 161280 0 161336 400
rect 162064 0 162120 400
rect 162848 0 162904 400
rect 163632 0 163688 400
rect 164416 0 164472 400
rect 165200 0 165256 400
rect 165984 0 166040 400
rect 166768 0 166824 400
rect 167552 0 167608 400
rect 168336 0 168392 400
rect 169120 0 169176 400
rect 169904 0 169960 400
rect 170688 0 170744 400
rect 171472 0 171528 400
rect 172256 0 172312 400
rect 173040 0 173096 400
rect 173824 0 173880 400
rect 174608 0 174664 400
rect 175392 0 175448 400
rect 176176 0 176232 400
rect 176960 0 177016 400
rect 177744 0 177800 400
rect 178528 0 178584 400
rect 179312 0 179368 400
rect 180096 0 180152 400
rect 180880 0 180936 400
rect 181664 0 181720 400
rect 182448 0 182504 400
rect 183232 0 183288 400
rect 184016 0 184072 400
rect 184800 0 184856 400
rect 185584 0 185640 400
rect 186368 0 186424 400
rect 187152 0 187208 400
rect 187936 0 187992 400
rect 188720 0 188776 400
rect 189504 0 189560 400
rect 190288 0 190344 400
rect 191072 0 191128 400
rect 191856 0 191912 400
rect 192640 0 192696 400
rect 193424 0 193480 400
rect 194208 0 194264 400
rect 194992 0 195048 400
rect 195776 0 195832 400
rect 196560 0 196616 400
rect 197344 0 197400 400
rect 198128 0 198184 400
rect 198912 0 198968 400
rect 199696 0 199752 400
rect 200480 0 200536 400
rect 201264 0 201320 400
rect 202048 0 202104 400
rect 202832 0 202888 400
rect 203616 0 203672 400
rect 204400 0 204456 400
rect 205184 0 205240 400
rect 205968 0 206024 400
rect 206752 0 206808 400
rect 207536 0 207592 400
rect 208320 0 208376 400
rect 209104 0 209160 400
rect 209888 0 209944 400
rect 210672 0 210728 400
rect 211456 0 211512 400
rect 212240 0 212296 400
rect 213024 0 213080 400
rect 213808 0 213864 400
rect 214592 0 214648 400
rect 215376 0 215432 400
rect 216160 0 216216 400
rect 216944 0 217000 400
rect 217728 0 217784 400
rect 218512 0 218568 400
rect 219296 0 219352 400
rect 220080 0 220136 400
rect 220864 0 220920 400
rect 221648 0 221704 400
rect 222432 0 222488 400
rect 223216 0 223272 400
rect 224000 0 224056 400
rect 224784 0 224840 400
rect 225568 0 225624 400
rect 226352 0 226408 400
rect 227136 0 227192 400
rect 227920 0 227976 400
rect 228704 0 228760 400
rect 229488 0 229544 400
rect 230272 0 230328 400
rect 231056 0 231112 400
rect 231840 0 231896 400
rect 232624 0 232680 400
rect 233408 0 233464 400
rect 234192 0 234248 400
rect 234976 0 235032 400
rect 235760 0 235816 400
rect 236544 0 236600 400
rect 237328 0 237384 400
rect 238112 0 238168 400
rect 238896 0 238952 400
rect 239680 0 239736 400
rect 240464 0 240520 400
rect 241248 0 241304 400
rect 242032 0 242088 400
rect 242816 0 242872 400
rect 243600 0 243656 400
rect 244384 0 244440 400
rect 245168 0 245224 400
rect 245952 0 246008 400
rect 246736 0 246792 400
rect 247520 0 247576 400
<< obsm2 >>
rect 966 430 258986 278339
rect 966 350 12290 430
rect 12406 350 13074 430
rect 13190 350 13858 430
rect 13974 350 14642 430
rect 14758 350 15426 430
rect 15542 350 16210 430
rect 16326 350 16994 430
rect 17110 350 17778 430
rect 17894 350 18562 430
rect 18678 350 19346 430
rect 19462 350 20130 430
rect 20246 350 20914 430
rect 21030 350 21698 430
rect 21814 350 22482 430
rect 22598 350 23266 430
rect 23382 350 24050 430
rect 24166 350 24834 430
rect 24950 350 25618 430
rect 25734 350 26402 430
rect 26518 350 27186 430
rect 27302 350 27970 430
rect 28086 350 28754 430
rect 28870 350 29538 430
rect 29654 350 30322 430
rect 30438 350 31106 430
rect 31222 350 31890 430
rect 32006 350 32674 430
rect 32790 350 33458 430
rect 33574 350 34242 430
rect 34358 350 35026 430
rect 35142 350 35810 430
rect 35926 350 36594 430
rect 36710 350 37378 430
rect 37494 350 38162 430
rect 38278 350 38946 430
rect 39062 350 39730 430
rect 39846 350 40514 430
rect 40630 350 41298 430
rect 41414 350 42082 430
rect 42198 350 42866 430
rect 42982 350 43650 430
rect 43766 350 44434 430
rect 44550 350 45218 430
rect 45334 350 46002 430
rect 46118 350 46786 430
rect 46902 350 47570 430
rect 47686 350 48354 430
rect 48470 350 49138 430
rect 49254 350 49922 430
rect 50038 350 50706 430
rect 50822 350 51490 430
rect 51606 350 52274 430
rect 52390 350 53058 430
rect 53174 350 53842 430
rect 53958 350 54626 430
rect 54742 350 55410 430
rect 55526 350 56194 430
rect 56310 350 56978 430
rect 57094 350 57762 430
rect 57878 350 58546 430
rect 58662 350 59330 430
rect 59446 350 60114 430
rect 60230 350 60898 430
rect 61014 350 61682 430
rect 61798 350 62466 430
rect 62582 350 63250 430
rect 63366 350 64034 430
rect 64150 350 64818 430
rect 64934 350 65602 430
rect 65718 350 66386 430
rect 66502 350 67170 430
rect 67286 350 67954 430
rect 68070 350 68738 430
rect 68854 350 69522 430
rect 69638 350 70306 430
rect 70422 350 71090 430
rect 71206 350 71874 430
rect 71990 350 72658 430
rect 72774 350 73442 430
rect 73558 350 74226 430
rect 74342 350 75010 430
rect 75126 350 75794 430
rect 75910 350 76578 430
rect 76694 350 77362 430
rect 77478 350 78146 430
rect 78262 350 78930 430
rect 79046 350 79714 430
rect 79830 350 80498 430
rect 80614 350 81282 430
rect 81398 350 82066 430
rect 82182 350 82850 430
rect 82966 350 83634 430
rect 83750 350 84418 430
rect 84534 350 85202 430
rect 85318 350 85986 430
rect 86102 350 86770 430
rect 86886 350 87554 430
rect 87670 350 88338 430
rect 88454 350 89122 430
rect 89238 350 89906 430
rect 90022 350 90690 430
rect 90806 350 91474 430
rect 91590 350 92258 430
rect 92374 350 93042 430
rect 93158 350 93826 430
rect 93942 350 94610 430
rect 94726 350 95394 430
rect 95510 350 96178 430
rect 96294 350 96962 430
rect 97078 350 97746 430
rect 97862 350 98530 430
rect 98646 350 99314 430
rect 99430 350 100098 430
rect 100214 350 100882 430
rect 100998 350 101666 430
rect 101782 350 102450 430
rect 102566 350 103234 430
rect 103350 350 104018 430
rect 104134 350 104802 430
rect 104918 350 105586 430
rect 105702 350 106370 430
rect 106486 350 107154 430
rect 107270 350 107938 430
rect 108054 350 108722 430
rect 108838 350 109506 430
rect 109622 350 110290 430
rect 110406 350 111074 430
rect 111190 350 111858 430
rect 111974 350 112642 430
rect 112758 350 113426 430
rect 113542 350 114210 430
rect 114326 350 114994 430
rect 115110 350 115778 430
rect 115894 350 116562 430
rect 116678 350 117346 430
rect 117462 350 118130 430
rect 118246 350 118914 430
rect 119030 350 119698 430
rect 119814 350 120482 430
rect 120598 350 121266 430
rect 121382 350 122050 430
rect 122166 350 122834 430
rect 122950 350 123618 430
rect 123734 350 124402 430
rect 124518 350 125186 430
rect 125302 350 125970 430
rect 126086 350 126754 430
rect 126870 350 127538 430
rect 127654 350 128322 430
rect 128438 350 129106 430
rect 129222 350 129890 430
rect 130006 350 130674 430
rect 130790 350 131458 430
rect 131574 350 132242 430
rect 132358 350 133026 430
rect 133142 350 133810 430
rect 133926 350 134594 430
rect 134710 350 135378 430
rect 135494 350 136162 430
rect 136278 350 136946 430
rect 137062 350 137730 430
rect 137846 350 138514 430
rect 138630 350 139298 430
rect 139414 350 140082 430
rect 140198 350 140866 430
rect 140982 350 141650 430
rect 141766 350 142434 430
rect 142550 350 143218 430
rect 143334 350 144002 430
rect 144118 350 144786 430
rect 144902 350 145570 430
rect 145686 350 146354 430
rect 146470 350 147138 430
rect 147254 350 147922 430
rect 148038 350 148706 430
rect 148822 350 149490 430
rect 149606 350 150274 430
rect 150390 350 151058 430
rect 151174 350 151842 430
rect 151958 350 152626 430
rect 152742 350 153410 430
rect 153526 350 154194 430
rect 154310 350 154978 430
rect 155094 350 155762 430
rect 155878 350 156546 430
rect 156662 350 157330 430
rect 157446 350 158114 430
rect 158230 350 158898 430
rect 159014 350 159682 430
rect 159798 350 160466 430
rect 160582 350 161250 430
rect 161366 350 162034 430
rect 162150 350 162818 430
rect 162934 350 163602 430
rect 163718 350 164386 430
rect 164502 350 165170 430
rect 165286 350 165954 430
rect 166070 350 166738 430
rect 166854 350 167522 430
rect 167638 350 168306 430
rect 168422 350 169090 430
rect 169206 350 169874 430
rect 169990 350 170658 430
rect 170774 350 171442 430
rect 171558 350 172226 430
rect 172342 350 173010 430
rect 173126 350 173794 430
rect 173910 350 174578 430
rect 174694 350 175362 430
rect 175478 350 176146 430
rect 176262 350 176930 430
rect 177046 350 177714 430
rect 177830 350 178498 430
rect 178614 350 179282 430
rect 179398 350 180066 430
rect 180182 350 180850 430
rect 180966 350 181634 430
rect 181750 350 182418 430
rect 182534 350 183202 430
rect 183318 350 183986 430
rect 184102 350 184770 430
rect 184886 350 185554 430
rect 185670 350 186338 430
rect 186454 350 187122 430
rect 187238 350 187906 430
rect 188022 350 188690 430
rect 188806 350 189474 430
rect 189590 350 190258 430
rect 190374 350 191042 430
rect 191158 350 191826 430
rect 191942 350 192610 430
rect 192726 350 193394 430
rect 193510 350 194178 430
rect 194294 350 194962 430
rect 195078 350 195746 430
rect 195862 350 196530 430
rect 196646 350 197314 430
rect 197430 350 198098 430
rect 198214 350 198882 430
rect 198998 350 199666 430
rect 199782 350 200450 430
rect 200566 350 201234 430
rect 201350 350 202018 430
rect 202134 350 202802 430
rect 202918 350 203586 430
rect 203702 350 204370 430
rect 204486 350 205154 430
rect 205270 350 205938 430
rect 206054 350 206722 430
rect 206838 350 207506 430
rect 207622 350 208290 430
rect 208406 350 209074 430
rect 209190 350 209858 430
rect 209974 350 210642 430
rect 210758 350 211426 430
rect 211542 350 212210 430
rect 212326 350 212994 430
rect 213110 350 213778 430
rect 213894 350 214562 430
rect 214678 350 215346 430
rect 215462 350 216130 430
rect 216246 350 216914 430
rect 217030 350 217698 430
rect 217814 350 218482 430
rect 218598 350 219266 430
rect 219382 350 220050 430
rect 220166 350 220834 430
rect 220950 350 221618 430
rect 221734 350 222402 430
rect 222518 350 223186 430
rect 223302 350 223970 430
rect 224086 350 224754 430
rect 224870 350 225538 430
rect 225654 350 226322 430
rect 226438 350 227106 430
rect 227222 350 227890 430
rect 228006 350 228674 430
rect 228790 350 229458 430
rect 229574 350 230242 430
rect 230358 350 231026 430
rect 231142 350 231810 430
rect 231926 350 232594 430
rect 232710 350 233378 430
rect 233494 350 234162 430
rect 234278 350 234946 430
rect 235062 350 235730 430
rect 235846 350 236514 430
rect 236630 350 237298 430
rect 237414 350 238082 430
rect 238198 350 238866 430
rect 238982 350 239650 430
rect 239766 350 240434 430
rect 240550 350 241218 430
rect 241334 350 242002 430
rect 242118 350 242786 430
rect 242902 350 243570 430
rect 243686 350 244354 430
rect 244470 350 245138 430
rect 245254 350 245922 430
rect 246038 350 246706 430
rect 246822 350 247490 430
rect 247606 350 258986 430
<< metal3 >>
rect 0 273840 400 273896
rect 259600 273840 260000 273896
rect 0 262192 400 262248
rect 259600 262192 260000 262248
rect 0 250544 400 250600
rect 259600 250544 260000 250600
rect 0 238896 400 238952
rect 259600 238896 260000 238952
rect 0 227248 400 227304
rect 259600 227248 260000 227304
rect 0 215600 400 215656
rect 259600 215600 260000 215656
rect 0 203952 400 204008
rect 259600 203952 260000 204008
rect 0 192304 400 192360
rect 259600 192304 260000 192360
rect 0 180656 400 180712
rect 259600 180656 260000 180712
rect 0 169008 400 169064
rect 259600 169008 260000 169064
rect 0 157360 400 157416
rect 259600 157360 260000 157416
rect 0 145712 400 145768
rect 259600 145712 260000 145768
rect 0 134064 400 134120
rect 259600 134064 260000 134120
rect 0 122416 400 122472
rect 259600 122416 260000 122472
rect 0 110768 400 110824
rect 259600 110768 260000 110824
rect 0 99120 400 99176
rect 259600 99120 260000 99176
rect 0 87472 400 87528
rect 259600 87472 260000 87528
rect 0 75824 400 75880
rect 259600 75824 260000 75880
rect 0 64176 400 64232
rect 259600 64176 260000 64232
rect 0 52528 400 52584
rect 259600 52528 260000 52584
rect 0 40880 400 40936
rect 259600 40880 260000 40936
rect 0 29232 400 29288
rect 259600 29232 260000 29288
rect 0 17584 400 17640
rect 259600 17584 260000 17640
rect 0 5936 400 5992
rect 259600 5936 260000 5992
<< obsm3 >>
rect 400 273926 259600 278334
rect 430 273810 259570 273926
rect 400 262278 259600 273810
rect 430 262162 259570 262278
rect 400 250630 259600 262162
rect 430 250514 259570 250630
rect 400 238982 259600 250514
rect 430 238866 259570 238982
rect 400 227334 259600 238866
rect 430 227218 259570 227334
rect 400 215686 259600 227218
rect 430 215570 259570 215686
rect 400 204038 259600 215570
rect 430 203922 259570 204038
rect 400 192390 259600 203922
rect 430 192274 259570 192390
rect 400 180742 259600 192274
rect 430 180626 259570 180742
rect 400 169094 259600 180626
rect 430 168978 259570 169094
rect 400 157446 259600 168978
rect 430 157330 259570 157446
rect 400 145798 259600 157330
rect 430 145682 259570 145798
rect 400 134150 259600 145682
rect 430 134034 259570 134150
rect 400 122502 259600 134034
rect 430 122386 259570 122502
rect 400 110854 259600 122386
rect 430 110738 259570 110854
rect 400 99206 259600 110738
rect 430 99090 259570 99206
rect 400 87558 259600 99090
rect 430 87442 259570 87558
rect 400 75910 259600 87442
rect 430 75794 259570 75910
rect 400 64262 259600 75794
rect 430 64146 259570 64262
rect 400 52614 259600 64146
rect 430 52498 259570 52614
rect 400 40966 259600 52498
rect 430 40850 259570 40966
rect 400 29318 259600 40850
rect 430 29202 259570 29318
rect 400 17670 259600 29202
rect 430 17554 259570 17670
rect 400 6022 259600 17554
rect 430 5906 259570 6022
rect 400 462 259600 5906
<< metal4 >>
rect 2224 1538 2384 278350
rect 9904 1538 10064 278350
rect 17584 1538 17744 278350
rect 25264 1538 25424 278350
rect 32944 1538 33104 278350
rect 40624 1538 40784 278350
rect 48304 1538 48464 278350
rect 55984 1538 56144 278350
rect 63664 1538 63824 278350
rect 71344 1538 71504 278350
rect 79024 1538 79184 278350
rect 86704 1538 86864 278350
rect 94384 1538 94544 278350
rect 102064 1538 102224 278350
rect 109744 1538 109904 278350
rect 117424 1538 117584 278350
rect 125104 1538 125264 278350
rect 132784 1538 132944 278350
rect 140464 1538 140624 278350
rect 148144 1538 148304 278350
rect 155824 1538 155984 278350
rect 163504 1538 163664 278350
rect 171184 1538 171344 278350
rect 178864 1538 179024 278350
rect 186544 1538 186704 278350
rect 194224 1538 194384 278350
rect 201904 1538 202064 278350
rect 209584 1538 209744 278350
rect 217264 1538 217424 278350
rect 224944 1538 225104 278350
rect 232624 1538 232784 278350
rect 240304 1538 240464 278350
rect 247984 1538 248144 278350
rect 255664 1538 255824 278350
<< obsm4 >>
rect 121758 2809 125074 4191
rect 125294 2809 132754 4191
rect 132974 2809 140434 4191
rect 140654 2809 148114 4191
rect 148334 2809 155794 4191
rect 156014 2809 162834 4191
<< labels >>
rlabel metal3 s 259600 5936 260000 5992 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 203952 400 204008 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 169008 400 169064 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 134064 400 134120 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 99120 400 99176 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 64176 400 64232 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 29232 400 29288 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 259600 40880 260000 40936 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 259600 75824 260000 75880 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 259600 110768 260000 110824 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 259600 145712 260000 145768 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 259600 180656 260000 180712 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 259600 215600 260000 215656 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 259600 250544 260000 250600 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 273840 400 273896 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 238896 400 238952 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 259600 29232 260000 29288 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 180656 400 180712 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 145712 400 145768 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 110768 400 110824 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 75824 400 75880 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 40880 400 40936 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 5936 400 5992 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 259600 64176 260000 64232 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 259600 99120 260000 99176 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 259600 134064 260000 134120 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 259600 169008 260000 169064 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 259600 203952 260000 204008 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 259600 238896 260000 238952 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 259600 273840 260000 273896 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 250544 400 250600 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 215600 400 215656 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 259600 17584 260000 17640 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 192304 400 192360 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 157360 400 157416 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 122416 400 122472 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 87472 400 87528 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 52528 400 52584 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 17584 400 17640 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 259600 52528 260000 52584 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 259600 87472 260000 87528 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 259600 122416 260000 122472 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 259600 157360 260000 157416 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 259600 192304 260000 192360 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 259600 227248 260000 227304 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 259600 262192 260000 262248 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 262192 400 262248 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 227248 400 227304 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 245952 0 246008 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 246736 0 246792 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 247520 0 247576 400 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 95424 0 95480 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 118944 0 119000 400 6 la_data_in[10]
port 53 nsew signal input
rlabel metal2 s 121296 0 121352 400 6 la_data_in[11]
port 54 nsew signal input
rlabel metal2 s 123648 0 123704 400 6 la_data_in[12]
port 55 nsew signal input
rlabel metal2 s 126000 0 126056 400 6 la_data_in[13]
port 56 nsew signal input
rlabel metal2 s 128352 0 128408 400 6 la_data_in[14]
port 57 nsew signal input
rlabel metal2 s 130704 0 130760 400 6 la_data_in[15]
port 58 nsew signal input
rlabel metal2 s 133056 0 133112 400 6 la_data_in[16]
port 59 nsew signal input
rlabel metal2 s 135408 0 135464 400 6 la_data_in[17]
port 60 nsew signal input
rlabel metal2 s 137760 0 137816 400 6 la_data_in[18]
port 61 nsew signal input
rlabel metal2 s 140112 0 140168 400 6 la_data_in[19]
port 62 nsew signal input
rlabel metal2 s 97776 0 97832 400 6 la_data_in[1]
port 63 nsew signal input
rlabel metal2 s 142464 0 142520 400 6 la_data_in[20]
port 64 nsew signal input
rlabel metal2 s 144816 0 144872 400 6 la_data_in[21]
port 65 nsew signal input
rlabel metal2 s 147168 0 147224 400 6 la_data_in[22]
port 66 nsew signal input
rlabel metal2 s 149520 0 149576 400 6 la_data_in[23]
port 67 nsew signal input
rlabel metal2 s 151872 0 151928 400 6 la_data_in[24]
port 68 nsew signal input
rlabel metal2 s 154224 0 154280 400 6 la_data_in[25]
port 69 nsew signal input
rlabel metal2 s 156576 0 156632 400 6 la_data_in[26]
port 70 nsew signal input
rlabel metal2 s 158928 0 158984 400 6 la_data_in[27]
port 71 nsew signal input
rlabel metal2 s 161280 0 161336 400 6 la_data_in[28]
port 72 nsew signal input
rlabel metal2 s 163632 0 163688 400 6 la_data_in[29]
port 73 nsew signal input
rlabel metal2 s 100128 0 100184 400 6 la_data_in[2]
port 74 nsew signal input
rlabel metal2 s 165984 0 166040 400 6 la_data_in[30]
port 75 nsew signal input
rlabel metal2 s 168336 0 168392 400 6 la_data_in[31]
port 76 nsew signal input
rlabel metal2 s 170688 0 170744 400 6 la_data_in[32]
port 77 nsew signal input
rlabel metal2 s 173040 0 173096 400 6 la_data_in[33]
port 78 nsew signal input
rlabel metal2 s 175392 0 175448 400 6 la_data_in[34]
port 79 nsew signal input
rlabel metal2 s 177744 0 177800 400 6 la_data_in[35]
port 80 nsew signal input
rlabel metal2 s 180096 0 180152 400 6 la_data_in[36]
port 81 nsew signal input
rlabel metal2 s 182448 0 182504 400 6 la_data_in[37]
port 82 nsew signal input
rlabel metal2 s 184800 0 184856 400 6 la_data_in[38]
port 83 nsew signal input
rlabel metal2 s 187152 0 187208 400 6 la_data_in[39]
port 84 nsew signal input
rlabel metal2 s 102480 0 102536 400 6 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 189504 0 189560 400 6 la_data_in[40]
port 86 nsew signal input
rlabel metal2 s 191856 0 191912 400 6 la_data_in[41]
port 87 nsew signal input
rlabel metal2 s 194208 0 194264 400 6 la_data_in[42]
port 88 nsew signal input
rlabel metal2 s 196560 0 196616 400 6 la_data_in[43]
port 89 nsew signal input
rlabel metal2 s 198912 0 198968 400 6 la_data_in[44]
port 90 nsew signal input
rlabel metal2 s 201264 0 201320 400 6 la_data_in[45]
port 91 nsew signal input
rlabel metal2 s 203616 0 203672 400 6 la_data_in[46]
port 92 nsew signal input
rlabel metal2 s 205968 0 206024 400 6 la_data_in[47]
port 93 nsew signal input
rlabel metal2 s 208320 0 208376 400 6 la_data_in[48]
port 94 nsew signal input
rlabel metal2 s 210672 0 210728 400 6 la_data_in[49]
port 95 nsew signal input
rlabel metal2 s 104832 0 104888 400 6 la_data_in[4]
port 96 nsew signal input
rlabel metal2 s 213024 0 213080 400 6 la_data_in[50]
port 97 nsew signal input
rlabel metal2 s 215376 0 215432 400 6 la_data_in[51]
port 98 nsew signal input
rlabel metal2 s 217728 0 217784 400 6 la_data_in[52]
port 99 nsew signal input
rlabel metal2 s 220080 0 220136 400 6 la_data_in[53]
port 100 nsew signal input
rlabel metal2 s 222432 0 222488 400 6 la_data_in[54]
port 101 nsew signal input
rlabel metal2 s 224784 0 224840 400 6 la_data_in[55]
port 102 nsew signal input
rlabel metal2 s 227136 0 227192 400 6 la_data_in[56]
port 103 nsew signal input
rlabel metal2 s 229488 0 229544 400 6 la_data_in[57]
port 104 nsew signal input
rlabel metal2 s 231840 0 231896 400 6 la_data_in[58]
port 105 nsew signal input
rlabel metal2 s 234192 0 234248 400 6 la_data_in[59]
port 106 nsew signal input
rlabel metal2 s 107184 0 107240 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 236544 0 236600 400 6 la_data_in[60]
port 108 nsew signal input
rlabel metal2 s 238896 0 238952 400 6 la_data_in[61]
port 109 nsew signal input
rlabel metal2 s 241248 0 241304 400 6 la_data_in[62]
port 110 nsew signal input
rlabel metal2 s 243600 0 243656 400 6 la_data_in[63]
port 111 nsew signal input
rlabel metal2 s 109536 0 109592 400 6 la_data_in[6]
port 112 nsew signal input
rlabel metal2 s 111888 0 111944 400 6 la_data_in[7]
port 113 nsew signal input
rlabel metal2 s 114240 0 114296 400 6 la_data_in[8]
port 114 nsew signal input
rlabel metal2 s 116592 0 116648 400 6 la_data_in[9]
port 115 nsew signal input
rlabel metal2 s 96208 0 96264 400 6 la_data_out[0]
port 116 nsew signal output
rlabel metal2 s 119728 0 119784 400 6 la_data_out[10]
port 117 nsew signal output
rlabel metal2 s 122080 0 122136 400 6 la_data_out[11]
port 118 nsew signal output
rlabel metal2 s 124432 0 124488 400 6 la_data_out[12]
port 119 nsew signal output
rlabel metal2 s 126784 0 126840 400 6 la_data_out[13]
port 120 nsew signal output
rlabel metal2 s 129136 0 129192 400 6 la_data_out[14]
port 121 nsew signal output
rlabel metal2 s 131488 0 131544 400 6 la_data_out[15]
port 122 nsew signal output
rlabel metal2 s 133840 0 133896 400 6 la_data_out[16]
port 123 nsew signal output
rlabel metal2 s 136192 0 136248 400 6 la_data_out[17]
port 124 nsew signal output
rlabel metal2 s 138544 0 138600 400 6 la_data_out[18]
port 125 nsew signal output
rlabel metal2 s 140896 0 140952 400 6 la_data_out[19]
port 126 nsew signal output
rlabel metal2 s 98560 0 98616 400 6 la_data_out[1]
port 127 nsew signal output
rlabel metal2 s 143248 0 143304 400 6 la_data_out[20]
port 128 nsew signal output
rlabel metal2 s 145600 0 145656 400 6 la_data_out[21]
port 129 nsew signal output
rlabel metal2 s 147952 0 148008 400 6 la_data_out[22]
port 130 nsew signal output
rlabel metal2 s 150304 0 150360 400 6 la_data_out[23]
port 131 nsew signal output
rlabel metal2 s 152656 0 152712 400 6 la_data_out[24]
port 132 nsew signal output
rlabel metal2 s 155008 0 155064 400 6 la_data_out[25]
port 133 nsew signal output
rlabel metal2 s 157360 0 157416 400 6 la_data_out[26]
port 134 nsew signal output
rlabel metal2 s 159712 0 159768 400 6 la_data_out[27]
port 135 nsew signal output
rlabel metal2 s 162064 0 162120 400 6 la_data_out[28]
port 136 nsew signal output
rlabel metal2 s 164416 0 164472 400 6 la_data_out[29]
port 137 nsew signal output
rlabel metal2 s 100912 0 100968 400 6 la_data_out[2]
port 138 nsew signal output
rlabel metal2 s 166768 0 166824 400 6 la_data_out[30]
port 139 nsew signal output
rlabel metal2 s 169120 0 169176 400 6 la_data_out[31]
port 140 nsew signal output
rlabel metal2 s 171472 0 171528 400 6 la_data_out[32]
port 141 nsew signal output
rlabel metal2 s 173824 0 173880 400 6 la_data_out[33]
port 142 nsew signal output
rlabel metal2 s 176176 0 176232 400 6 la_data_out[34]
port 143 nsew signal output
rlabel metal2 s 178528 0 178584 400 6 la_data_out[35]
port 144 nsew signal output
rlabel metal2 s 180880 0 180936 400 6 la_data_out[36]
port 145 nsew signal output
rlabel metal2 s 183232 0 183288 400 6 la_data_out[37]
port 146 nsew signal output
rlabel metal2 s 185584 0 185640 400 6 la_data_out[38]
port 147 nsew signal output
rlabel metal2 s 187936 0 187992 400 6 la_data_out[39]
port 148 nsew signal output
rlabel metal2 s 103264 0 103320 400 6 la_data_out[3]
port 149 nsew signal output
rlabel metal2 s 190288 0 190344 400 6 la_data_out[40]
port 150 nsew signal output
rlabel metal2 s 192640 0 192696 400 6 la_data_out[41]
port 151 nsew signal output
rlabel metal2 s 194992 0 195048 400 6 la_data_out[42]
port 152 nsew signal output
rlabel metal2 s 197344 0 197400 400 6 la_data_out[43]
port 153 nsew signal output
rlabel metal2 s 199696 0 199752 400 6 la_data_out[44]
port 154 nsew signal output
rlabel metal2 s 202048 0 202104 400 6 la_data_out[45]
port 155 nsew signal output
rlabel metal2 s 204400 0 204456 400 6 la_data_out[46]
port 156 nsew signal output
rlabel metal2 s 206752 0 206808 400 6 la_data_out[47]
port 157 nsew signal output
rlabel metal2 s 209104 0 209160 400 6 la_data_out[48]
port 158 nsew signal output
rlabel metal2 s 211456 0 211512 400 6 la_data_out[49]
port 159 nsew signal output
rlabel metal2 s 105616 0 105672 400 6 la_data_out[4]
port 160 nsew signal output
rlabel metal2 s 213808 0 213864 400 6 la_data_out[50]
port 161 nsew signal output
rlabel metal2 s 216160 0 216216 400 6 la_data_out[51]
port 162 nsew signal output
rlabel metal2 s 218512 0 218568 400 6 la_data_out[52]
port 163 nsew signal output
rlabel metal2 s 220864 0 220920 400 6 la_data_out[53]
port 164 nsew signal output
rlabel metal2 s 223216 0 223272 400 6 la_data_out[54]
port 165 nsew signal output
rlabel metal2 s 225568 0 225624 400 6 la_data_out[55]
port 166 nsew signal output
rlabel metal2 s 227920 0 227976 400 6 la_data_out[56]
port 167 nsew signal output
rlabel metal2 s 230272 0 230328 400 6 la_data_out[57]
port 168 nsew signal output
rlabel metal2 s 232624 0 232680 400 6 la_data_out[58]
port 169 nsew signal output
rlabel metal2 s 234976 0 235032 400 6 la_data_out[59]
port 170 nsew signal output
rlabel metal2 s 107968 0 108024 400 6 la_data_out[5]
port 171 nsew signal output
rlabel metal2 s 237328 0 237384 400 6 la_data_out[60]
port 172 nsew signal output
rlabel metal2 s 239680 0 239736 400 6 la_data_out[61]
port 173 nsew signal output
rlabel metal2 s 242032 0 242088 400 6 la_data_out[62]
port 174 nsew signal output
rlabel metal2 s 244384 0 244440 400 6 la_data_out[63]
port 175 nsew signal output
rlabel metal2 s 110320 0 110376 400 6 la_data_out[6]
port 176 nsew signal output
rlabel metal2 s 112672 0 112728 400 6 la_data_out[7]
port 177 nsew signal output
rlabel metal2 s 115024 0 115080 400 6 la_data_out[8]
port 178 nsew signal output
rlabel metal2 s 117376 0 117432 400 6 la_data_out[9]
port 179 nsew signal output
rlabel metal2 s 96992 0 97048 400 6 la_oenb[0]
port 180 nsew signal input
rlabel metal2 s 120512 0 120568 400 6 la_oenb[10]
port 181 nsew signal input
rlabel metal2 s 122864 0 122920 400 6 la_oenb[11]
port 182 nsew signal input
rlabel metal2 s 125216 0 125272 400 6 la_oenb[12]
port 183 nsew signal input
rlabel metal2 s 127568 0 127624 400 6 la_oenb[13]
port 184 nsew signal input
rlabel metal2 s 129920 0 129976 400 6 la_oenb[14]
port 185 nsew signal input
rlabel metal2 s 132272 0 132328 400 6 la_oenb[15]
port 186 nsew signal input
rlabel metal2 s 134624 0 134680 400 6 la_oenb[16]
port 187 nsew signal input
rlabel metal2 s 136976 0 137032 400 6 la_oenb[17]
port 188 nsew signal input
rlabel metal2 s 139328 0 139384 400 6 la_oenb[18]
port 189 nsew signal input
rlabel metal2 s 141680 0 141736 400 6 la_oenb[19]
port 190 nsew signal input
rlabel metal2 s 99344 0 99400 400 6 la_oenb[1]
port 191 nsew signal input
rlabel metal2 s 144032 0 144088 400 6 la_oenb[20]
port 192 nsew signal input
rlabel metal2 s 146384 0 146440 400 6 la_oenb[21]
port 193 nsew signal input
rlabel metal2 s 148736 0 148792 400 6 la_oenb[22]
port 194 nsew signal input
rlabel metal2 s 151088 0 151144 400 6 la_oenb[23]
port 195 nsew signal input
rlabel metal2 s 153440 0 153496 400 6 la_oenb[24]
port 196 nsew signal input
rlabel metal2 s 155792 0 155848 400 6 la_oenb[25]
port 197 nsew signal input
rlabel metal2 s 158144 0 158200 400 6 la_oenb[26]
port 198 nsew signal input
rlabel metal2 s 160496 0 160552 400 6 la_oenb[27]
port 199 nsew signal input
rlabel metal2 s 162848 0 162904 400 6 la_oenb[28]
port 200 nsew signal input
rlabel metal2 s 165200 0 165256 400 6 la_oenb[29]
port 201 nsew signal input
rlabel metal2 s 101696 0 101752 400 6 la_oenb[2]
port 202 nsew signal input
rlabel metal2 s 167552 0 167608 400 6 la_oenb[30]
port 203 nsew signal input
rlabel metal2 s 169904 0 169960 400 6 la_oenb[31]
port 204 nsew signal input
rlabel metal2 s 172256 0 172312 400 6 la_oenb[32]
port 205 nsew signal input
rlabel metal2 s 174608 0 174664 400 6 la_oenb[33]
port 206 nsew signal input
rlabel metal2 s 176960 0 177016 400 6 la_oenb[34]
port 207 nsew signal input
rlabel metal2 s 179312 0 179368 400 6 la_oenb[35]
port 208 nsew signal input
rlabel metal2 s 181664 0 181720 400 6 la_oenb[36]
port 209 nsew signal input
rlabel metal2 s 184016 0 184072 400 6 la_oenb[37]
port 210 nsew signal input
rlabel metal2 s 186368 0 186424 400 6 la_oenb[38]
port 211 nsew signal input
rlabel metal2 s 188720 0 188776 400 6 la_oenb[39]
port 212 nsew signal input
rlabel metal2 s 104048 0 104104 400 6 la_oenb[3]
port 213 nsew signal input
rlabel metal2 s 191072 0 191128 400 6 la_oenb[40]
port 214 nsew signal input
rlabel metal2 s 193424 0 193480 400 6 la_oenb[41]
port 215 nsew signal input
rlabel metal2 s 195776 0 195832 400 6 la_oenb[42]
port 216 nsew signal input
rlabel metal2 s 198128 0 198184 400 6 la_oenb[43]
port 217 nsew signal input
rlabel metal2 s 200480 0 200536 400 6 la_oenb[44]
port 218 nsew signal input
rlabel metal2 s 202832 0 202888 400 6 la_oenb[45]
port 219 nsew signal input
rlabel metal2 s 205184 0 205240 400 6 la_oenb[46]
port 220 nsew signal input
rlabel metal2 s 207536 0 207592 400 6 la_oenb[47]
port 221 nsew signal input
rlabel metal2 s 209888 0 209944 400 6 la_oenb[48]
port 222 nsew signal input
rlabel metal2 s 212240 0 212296 400 6 la_oenb[49]
port 223 nsew signal input
rlabel metal2 s 106400 0 106456 400 6 la_oenb[4]
port 224 nsew signal input
rlabel metal2 s 214592 0 214648 400 6 la_oenb[50]
port 225 nsew signal input
rlabel metal2 s 216944 0 217000 400 6 la_oenb[51]
port 226 nsew signal input
rlabel metal2 s 219296 0 219352 400 6 la_oenb[52]
port 227 nsew signal input
rlabel metal2 s 221648 0 221704 400 6 la_oenb[53]
port 228 nsew signal input
rlabel metal2 s 224000 0 224056 400 6 la_oenb[54]
port 229 nsew signal input
rlabel metal2 s 226352 0 226408 400 6 la_oenb[55]
port 230 nsew signal input
rlabel metal2 s 228704 0 228760 400 6 la_oenb[56]
port 231 nsew signal input
rlabel metal2 s 231056 0 231112 400 6 la_oenb[57]
port 232 nsew signal input
rlabel metal2 s 233408 0 233464 400 6 la_oenb[58]
port 233 nsew signal input
rlabel metal2 s 235760 0 235816 400 6 la_oenb[59]
port 234 nsew signal input
rlabel metal2 s 108752 0 108808 400 6 la_oenb[5]
port 235 nsew signal input
rlabel metal2 s 238112 0 238168 400 6 la_oenb[60]
port 236 nsew signal input
rlabel metal2 s 240464 0 240520 400 6 la_oenb[61]
port 237 nsew signal input
rlabel metal2 s 242816 0 242872 400 6 la_oenb[62]
port 238 nsew signal input
rlabel metal2 s 245168 0 245224 400 6 la_oenb[63]
port 239 nsew signal input
rlabel metal2 s 111104 0 111160 400 6 la_oenb[6]
port 240 nsew signal input
rlabel metal2 s 113456 0 113512 400 6 la_oenb[7]
port 241 nsew signal input
rlabel metal2 s 115808 0 115864 400 6 la_oenb[8]
port 242 nsew signal input
rlabel metal2 s 118160 0 118216 400 6 la_oenb[9]
port 243 nsew signal input
rlabel metal4 s 2224 1538 2384 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 278350 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 278350 6 vss
port 245 nsew ground bidirectional
rlabel metal2 s 12320 0 12376 400 6 wb_clk_i
port 246 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 wb_rst_i
port 247 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 wbs_ack_o
port 248 nsew signal output
rlabel metal2 s 17024 0 17080 400 6 wbs_adr_i[0]
port 249 nsew signal input
rlabel metal2 s 43680 0 43736 400 6 wbs_adr_i[10]
port 250 nsew signal input
rlabel metal2 s 46032 0 46088 400 6 wbs_adr_i[11]
port 251 nsew signal input
rlabel metal2 s 48384 0 48440 400 6 wbs_adr_i[12]
port 252 nsew signal input
rlabel metal2 s 50736 0 50792 400 6 wbs_adr_i[13]
port 253 nsew signal input
rlabel metal2 s 53088 0 53144 400 6 wbs_adr_i[14]
port 254 nsew signal input
rlabel metal2 s 55440 0 55496 400 6 wbs_adr_i[15]
port 255 nsew signal input
rlabel metal2 s 57792 0 57848 400 6 wbs_adr_i[16]
port 256 nsew signal input
rlabel metal2 s 60144 0 60200 400 6 wbs_adr_i[17]
port 257 nsew signal input
rlabel metal2 s 62496 0 62552 400 6 wbs_adr_i[18]
port 258 nsew signal input
rlabel metal2 s 64848 0 64904 400 6 wbs_adr_i[19]
port 259 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 wbs_adr_i[1]
port 260 nsew signal input
rlabel metal2 s 67200 0 67256 400 6 wbs_adr_i[20]
port 261 nsew signal input
rlabel metal2 s 69552 0 69608 400 6 wbs_adr_i[21]
port 262 nsew signal input
rlabel metal2 s 71904 0 71960 400 6 wbs_adr_i[22]
port 263 nsew signal input
rlabel metal2 s 74256 0 74312 400 6 wbs_adr_i[23]
port 264 nsew signal input
rlabel metal2 s 76608 0 76664 400 6 wbs_adr_i[24]
port 265 nsew signal input
rlabel metal2 s 78960 0 79016 400 6 wbs_adr_i[25]
port 266 nsew signal input
rlabel metal2 s 81312 0 81368 400 6 wbs_adr_i[26]
port 267 nsew signal input
rlabel metal2 s 83664 0 83720 400 6 wbs_adr_i[27]
port 268 nsew signal input
rlabel metal2 s 86016 0 86072 400 6 wbs_adr_i[28]
port 269 nsew signal input
rlabel metal2 s 88368 0 88424 400 6 wbs_adr_i[29]
port 270 nsew signal input
rlabel metal2 s 23296 0 23352 400 6 wbs_adr_i[2]
port 271 nsew signal input
rlabel metal2 s 90720 0 90776 400 6 wbs_adr_i[30]
port 272 nsew signal input
rlabel metal2 s 93072 0 93128 400 6 wbs_adr_i[31]
port 273 nsew signal input
rlabel metal2 s 26432 0 26488 400 6 wbs_adr_i[3]
port 274 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 wbs_adr_i[4]
port 275 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 wbs_adr_i[5]
port 276 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 wbs_adr_i[6]
port 277 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 wbs_adr_i[7]
port 278 nsew signal input
rlabel metal2 s 38976 0 39032 400 6 wbs_adr_i[8]
port 279 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 wbs_adr_i[9]
port 280 nsew signal input
rlabel metal2 s 14672 0 14728 400 6 wbs_cyc_i
port 281 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 wbs_dat_i[0]
port 282 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 wbs_dat_i[10]
port 283 nsew signal input
rlabel metal2 s 46816 0 46872 400 6 wbs_dat_i[11]
port 284 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 wbs_dat_i[12]
port 285 nsew signal input
rlabel metal2 s 51520 0 51576 400 6 wbs_dat_i[13]
port 286 nsew signal input
rlabel metal2 s 53872 0 53928 400 6 wbs_dat_i[14]
port 287 nsew signal input
rlabel metal2 s 56224 0 56280 400 6 wbs_dat_i[15]
port 288 nsew signal input
rlabel metal2 s 58576 0 58632 400 6 wbs_dat_i[16]
port 289 nsew signal input
rlabel metal2 s 60928 0 60984 400 6 wbs_dat_i[17]
port 290 nsew signal input
rlabel metal2 s 63280 0 63336 400 6 wbs_dat_i[18]
port 291 nsew signal input
rlabel metal2 s 65632 0 65688 400 6 wbs_dat_i[19]
port 292 nsew signal input
rlabel metal2 s 20944 0 21000 400 6 wbs_dat_i[1]
port 293 nsew signal input
rlabel metal2 s 67984 0 68040 400 6 wbs_dat_i[20]
port 294 nsew signal input
rlabel metal2 s 70336 0 70392 400 6 wbs_dat_i[21]
port 295 nsew signal input
rlabel metal2 s 72688 0 72744 400 6 wbs_dat_i[22]
port 296 nsew signal input
rlabel metal2 s 75040 0 75096 400 6 wbs_dat_i[23]
port 297 nsew signal input
rlabel metal2 s 77392 0 77448 400 6 wbs_dat_i[24]
port 298 nsew signal input
rlabel metal2 s 79744 0 79800 400 6 wbs_dat_i[25]
port 299 nsew signal input
rlabel metal2 s 82096 0 82152 400 6 wbs_dat_i[26]
port 300 nsew signal input
rlabel metal2 s 84448 0 84504 400 6 wbs_dat_i[27]
port 301 nsew signal input
rlabel metal2 s 86800 0 86856 400 6 wbs_dat_i[28]
port 302 nsew signal input
rlabel metal2 s 89152 0 89208 400 6 wbs_dat_i[29]
port 303 nsew signal input
rlabel metal2 s 24080 0 24136 400 6 wbs_dat_i[2]
port 304 nsew signal input
rlabel metal2 s 91504 0 91560 400 6 wbs_dat_i[30]
port 305 nsew signal input
rlabel metal2 s 93856 0 93912 400 6 wbs_dat_i[31]
port 306 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 wbs_dat_i[3]
port 307 nsew signal input
rlabel metal2 s 30352 0 30408 400 6 wbs_dat_i[4]
port 308 nsew signal input
rlabel metal2 s 32704 0 32760 400 6 wbs_dat_i[5]
port 309 nsew signal input
rlabel metal2 s 35056 0 35112 400 6 wbs_dat_i[6]
port 310 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 wbs_dat_i[7]
port 311 nsew signal input
rlabel metal2 s 39760 0 39816 400 6 wbs_dat_i[8]
port 312 nsew signal input
rlabel metal2 s 42112 0 42168 400 6 wbs_dat_i[9]
port 313 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 wbs_dat_o[0]
port 314 nsew signal output
rlabel metal2 s 45248 0 45304 400 6 wbs_dat_o[10]
port 315 nsew signal output
rlabel metal2 s 47600 0 47656 400 6 wbs_dat_o[11]
port 316 nsew signal output
rlabel metal2 s 49952 0 50008 400 6 wbs_dat_o[12]
port 317 nsew signal output
rlabel metal2 s 52304 0 52360 400 6 wbs_dat_o[13]
port 318 nsew signal output
rlabel metal2 s 54656 0 54712 400 6 wbs_dat_o[14]
port 319 nsew signal output
rlabel metal2 s 57008 0 57064 400 6 wbs_dat_o[15]
port 320 nsew signal output
rlabel metal2 s 59360 0 59416 400 6 wbs_dat_o[16]
port 321 nsew signal output
rlabel metal2 s 61712 0 61768 400 6 wbs_dat_o[17]
port 322 nsew signal output
rlabel metal2 s 64064 0 64120 400 6 wbs_dat_o[18]
port 323 nsew signal output
rlabel metal2 s 66416 0 66472 400 6 wbs_dat_o[19]
port 324 nsew signal output
rlabel metal2 s 21728 0 21784 400 6 wbs_dat_o[1]
port 325 nsew signal output
rlabel metal2 s 68768 0 68824 400 6 wbs_dat_o[20]
port 326 nsew signal output
rlabel metal2 s 71120 0 71176 400 6 wbs_dat_o[21]
port 327 nsew signal output
rlabel metal2 s 73472 0 73528 400 6 wbs_dat_o[22]
port 328 nsew signal output
rlabel metal2 s 75824 0 75880 400 6 wbs_dat_o[23]
port 329 nsew signal output
rlabel metal2 s 78176 0 78232 400 6 wbs_dat_o[24]
port 330 nsew signal output
rlabel metal2 s 80528 0 80584 400 6 wbs_dat_o[25]
port 331 nsew signal output
rlabel metal2 s 82880 0 82936 400 6 wbs_dat_o[26]
port 332 nsew signal output
rlabel metal2 s 85232 0 85288 400 6 wbs_dat_o[27]
port 333 nsew signal output
rlabel metal2 s 87584 0 87640 400 6 wbs_dat_o[28]
port 334 nsew signal output
rlabel metal2 s 89936 0 89992 400 6 wbs_dat_o[29]
port 335 nsew signal output
rlabel metal2 s 24864 0 24920 400 6 wbs_dat_o[2]
port 336 nsew signal output
rlabel metal2 s 92288 0 92344 400 6 wbs_dat_o[30]
port 337 nsew signal output
rlabel metal2 s 94640 0 94696 400 6 wbs_dat_o[31]
port 338 nsew signal output
rlabel metal2 s 28000 0 28056 400 6 wbs_dat_o[3]
port 339 nsew signal output
rlabel metal2 s 31136 0 31192 400 6 wbs_dat_o[4]
port 340 nsew signal output
rlabel metal2 s 33488 0 33544 400 6 wbs_dat_o[5]
port 341 nsew signal output
rlabel metal2 s 35840 0 35896 400 6 wbs_dat_o[6]
port 342 nsew signal output
rlabel metal2 s 38192 0 38248 400 6 wbs_dat_o[7]
port 343 nsew signal output
rlabel metal2 s 40544 0 40600 400 6 wbs_dat_o[8]
port 344 nsew signal output
rlabel metal2 s 42896 0 42952 400 6 wbs_dat_o[9]
port 345 nsew signal output
rlabel metal2 s 19376 0 19432 400 6 wbs_sel_i[0]
port 346 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 wbs_sel_i[1]
port 347 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 wbs_sel_i[2]
port 348 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_sel_i[3]
port 349 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 wbs_stb_i
port 350 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 wbs_we_i
port 351 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 260000 280000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23052858
string GDS_FILE /home/yatharth/gf180_project/caravel_user_project/openlane/user_proj_example/runs/23_12_04_11_57/results/signoff/user_proj_example.magic.gds
string GDS_START 280538
<< end >>

